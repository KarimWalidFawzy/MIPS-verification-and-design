
module MIPS();
    ALU alu(/*pins inserted*/);
endmodule