module Controlbits(
    input opcode[3:0]
);
    
endmodule