interface MIPSifc;
    
endinterface